module i8_trunc(
    input [11:0] A,
    output [3:0] B
);

endmodule

