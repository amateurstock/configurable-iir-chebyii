module i8_trunc(
    input [7:0] A,
    output [3:0] B
);

endmodule

