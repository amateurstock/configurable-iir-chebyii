module i36_delay(
);

endmodule

